`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:45:19 10/06/2017 
// Design Name: 
// Module Name:    ins_deco 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ins_deco(
    output wr_pc,
    output [1:0] sel_a,
    output sel_b,
    output wr_acc,
    output op,
    output wr_ram,
    output rd_ram,
    input [4:0] opcode
    );


endmodule
